library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity shift_rows is 
    port (
    i_state_in  : in std_ulogic_vector(127 downto 0);
    o_state_out : out std_ulogic_vector(127 downto 0)
    );
end entity shift_rows;
